module registers (
        input logic [4:0] read_register1, read_register2, write_register,
        input logic [31:0] write_data,
        input logic RegWrite,
        output logic [31:0] read_data1, read_data2
    );

    /** LÓGICA INTERNA DO REGISTRADOR **/

endmodule